module duplicate_name ();  
    wire unconnected_wire; // This wire is unconnected

endmodule

module duplicate_name ();  // Duplicate module name
    logic x;
endmodule