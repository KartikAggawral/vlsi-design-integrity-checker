module and_gate (
    input wire a,      // First input
    input wire b,      // Second input
    output wire out    // Output
);

    assign out = a & b;  // AND gate operation

endmodule
